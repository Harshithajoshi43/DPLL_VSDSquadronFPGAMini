  GNU nano 7.2                                                                                                      sim_lib.v                                                                                                                
// sim_lib.v — stub for the Lattice SB_GB primitive
module SB_GB (
    input  USER_SIGNAL_TO_GLOBAL_BUFFER,
    output GLOBAL_BUFFER_OUTPUT
);
  assign GLOBAL_BUFFER_OUTPUT = USER_SIGNAL_TO_GLOBAL_BUFFER;
endmodule
